

`timescale 1ns / 1ps
`default_nettype none


module tb_vdma_axi4_to_axi4s_core();
	
	
	parameter	RATE = 1000.0/50.0;
	
	reg		clk   = 1'b0;
	always #(RATE/2.0)	clk = ~clk;
	
	reg		reset = 1'b1;
	initial #(RATE*100)	reset <= 1'b0;
	
	
	initial begin
		$dumpfile("tb_vdma_axi4_to_axi4s_core.vcd");
		$dumpvars(0, tb_vdma_axi4_to_axi4s_core);
	#(RATE*640*480*3*2)
		$finish;
	end
	
	
	
	parameter	AXI4_ID_WIDTH    = 6;
	parameter	AXI4_ADDR_WIDTH  = 32;
	parameter	AXI4_LEN_WIDTH   = 8;
	parameter	AXI4_QOS_WIDTH   = 4;
	parameter	AXI4S_USER_WIDTH = 1;
	parameter	AXI4S_DATA_WIDTH = 24;
	parameter	STRIDE_WIDTH     = 12;
	parameter	INDEX_WIDTH      = 8;
	parameter	H_WIDTH          = 12;
	parameter	V_WIDTH          = 12;
	
	wire							enable = 1'b1;
	wire							busy;
	
	wire	[AXI4_ADDR_WIDTH-1:0]	param_addr   = 0;
	wire	[STRIDE_WIDTH-1:0]		param_stride = 4096;
	wire	[H_WIDTH-1:0]			param_width  = 640;
	wire	[V_WIDTH-1:0]			param_height = 480;
	wire	[AXI4_LEN_WIDTH-1:0]	param_arlen  = 7;
	
	wire	[INDEX_WIDTH-1:0]		status_index;
	wire	[AXI4_ADDR_WIDTH-1:0]	status_addr;
	wire	[STRIDE_WIDTH-1:0]		status_stride;
	wire	[H_WIDTH-1:0]			status_width;
	wire	[V_WIDTH-1:0]			status_height;
	wire	[AXI4_LEN_WIDTH-1:0]	status_arlen;
	
	wire	[AXI4_ID_WIDTH-1:0]		axi4_arid;
	wire	[AXI4_ADDR_WIDTH-1:0]	axi4_araddr;
	wire	[1:0]					axi4_arburst;
	wire	[3:0]					axi4_arcache;
	wire	[AXI4_LEN_WIDTH-1:0]	axi4_arlen;
	wire	[0:0]					axi4_arlock;
	wire	[2:0]					axi4_arprot;
	wire	[AXI4_QOS_WIDTH-1:0]	axi4_arqos;
	wire	[3:0]					axi4_arregion;
	wire	[2:0]					axi4_arsize;
	wire							axi4_arvalid;
	wire							axi4_arready;
	wire	[AXI4_ID_WIDTH-1:0]		axi4_rid;
	wire	[1:0]					axi4_rresp;
	wire	[31:0]					axi4_rdata;
	wire							axi4_rlast;
	wire							axi4_rvalid;
	wire							axi4_rready;
	
	wire	[AXI4S_USER_WIDTH-1:0]	axi4s_tuser;
	wire							axi4s_tlast;
	wire	[AXI4S_DATA_WIDTH-1:0]	axi4s_tdata;
	wire							axi4s_tvalid;
	wire							axi4s_tready = 1'b1;
	
	vdma_axi4_to_axi4s_core
			#(
				.AXI4_ID_WIDTH		(AXI4_ID_WIDTH),
				.AXI4_ADDR_WIDTH	(AXI4_ADDR_WIDTH),
				.AXI4_LEN_WIDTH		(AXI4_LEN_WIDTH),
				.AXI4_QOS_WIDTH		(AXI4_QOS_WIDTH),
				.AXI4S_USER_WIDTH	(AXI4S_USER_WIDTH),
				.AXI4S_DATA_WIDTH	(AXI4S_DATA_WIDTH),
				.STRIDE_WIDTH		(STRIDE_WIDTH),
				.INDEX_WIDTH		(INDEX_WIDTH),
				.H_WIDTH			(H_WIDTH),
				.V_WIDTH			(V_WIDTH)
			)
		i_vdma_axi4_to_axi4s_core
			(
				.aresetn			(~reset),
				.aclk				(clk),
				
				.ctl_enable			(enable),
				.ctl_update			(1'b1),
				.ctl_busy			(busy),
				.ctl_index			(status_index),
				
				.param_addr			(param_addr),
				.param_stride		(param_stride),
				.param_width		(param_width),
				.param_height		(param_height),
				.param_arlen		(param_arlen),
				
				.monitor_addr		(status_addr),
				.monitor_stride		(status_stride),
				.monitor_width		(status_width),
				.monitor_height		(status_height),
				.monitor_arlen		(status_arlen),
				
				.m_axi4_arid		(axi4_arid),
				.m_axi4_araddr		(axi4_araddr),
				.m_axi4_arburst		(axi4_arburst),
				.m_axi4_arcache		(axi4_arcache),
				.m_axi4_arlen		(axi4_arlen),
				.m_axi4_arlock		(axi4_arlock),
				.m_axi4_arprot		(axi4_arprot),
				.m_axi4_arqos		(axi4_arqos),
				.m_axi4_arregion	(axi4_arregion),
				.m_axi4_arsize		(axi4_arsize),
				.m_axi4_arvalid		(axi4_arvalid),
				.m_axi4_arready		(axi4_arready),
				.m_axi4_rid			(axi4_rid),
				.m_axi4_rresp		(axi4_rresp),
				.m_axi4_rdata		(axi4_rdata),
				.m_axi4_rlast		(axi4_rlast),
				.m_axi4_rvalid		(axi4_rvalid),
				.m_axi4_rready		(axi4_rready),
				
				.m_axi4s_tuser		(axi4s_tuser),
				.m_axi4s_tlast		(axi4s_tlast),
				.m_axi4s_tdata		(axi4s_tdata),
				.m_axi4s_tvalid		(axi4s_tvalid),
				.m_axi4s_tready		(axi4s_tready)
			);
	



	parameter	AXI4_DATA_SIZE   = 2;	// 0:8bit, 1:16bit, 2:32bit ...
	parameter	AXI4_DATA_WIDTH  = (8 << AXI4_DATA_SIZE);
	parameter	AXI4_STRB_WIDTH  = (1 << AXI4_DATA_SIZE);

	// master AXI4 (write)
	wire	[AXI4_ID_WIDTH-1:0]		axi4_awid;
	wire	[AXI4_ADDR_WIDTH-1:0]	axi4_awaddr;
	wire	[1:0]					axi4_awburst;
	wire	[3:0]					axi4_awcache;
	wire	[AXI4_LEN_WIDTH-1:0]	axi4_awlen;
	wire	[0:0]					axi4_awlock;
	wire	[2:0]					axi4_awprot;
	wire	[AXI4_QOS_WIDTH-1:0]	axi4_awqos;
	wire	[3:0]					axi4_awregion;
	wire	[2:0]					axi4_awsize;
	wire							axi4_awvalid;
	wire							axi4_awready;
	
	wire	[AXI4_STRB_WIDTH-1:0]	axi4_wstrb;
	wire	[AXI4_DATA_WIDTH-1:0]	axi4_wdata;
	wire							axi4_wlast;
	wire							axi4_wvalid;
	wire							axi4_wready;
	
	wire	[AXI4_ID_WIDTH-1:0]		axi4_bid;
	wire	[1:0]					axi4_bresp;
	wire							axi4_bvalid;
	wire							axi4_bready;
	
	// slave AXI4-Stream (output)
	wire	[AXI4S_USER_WIDTH-1:0]	s_axi4s_tuser;
	wire							s_axi4s_tlast;
	wire	[31:0]					s_axi4s_tdata;
	wire							s_axi4s_tvalid;
	wire							s_axi4s_tready;
	
	
	reg		[3:1]					rand;
	reg								s_axi4s_busy;
	always @(posedge clk) begin
		rand         <= $random;
		s_axi4s_busy <= (rand == 0);
	end
	
	model_axi4s_master
			#(
				.AXI4S_DATA_WIDTH	(32),
				.X_NUM				(640),
				.Y_NUM				(480)
			)
		i_model_axi4s_master
			(
				.aresetn			(~reset),
				.aclk				(clk),
				
				.m_axi4s_tuser		(s_axi4s_tuser),
				.m_axi4s_tlast		(s_axi4s_tlast),
				.m_axi4s_tdata		(s_axi4s_tdata),
				.m_axi4s_tvalid		(s_axi4s_tvalid),
				.m_axi4s_tready		(s_axi4s_tready & ~s_axi4s_busy)
			);
	
	
	vdma_axi4s_to_axi4_core
			#(
				.AXI4_ID_WIDTH		(AXI4_ID_WIDTH),
				.AXI4_ADDR_WIDTH	(AXI4_ADDR_WIDTH),
				.AXI4_LEN_WIDTH		(AXI4_LEN_WIDTH),
				.AXI4_QOS_WIDTH		(AXI4_QOS_WIDTH),
				.AXI4_DATA_SIZE		(AXI4_DATA_SIZE),
				.AXI4S_USER_WIDTH	(1),
				.AXI4S_DATA_WIDTH	(32),
				.STRIDE_WIDTH		(14),
				.INDEX_WIDTH		(8),
				.H_WIDTH			(12),
				.V_WIDTH			(12)
			)
		i_vdma_axi4s_to_axi4_core
			(
				.aresetn			(~reset),
				.aclk				(clk),
				
				.ctl_enable			(1'b1),
				.ctl_update			(1'b1),
				.ctl_busy			(),
				.ctl_index			(),
				
				.param_addr			(32'h0),
				.param_stride		(640),
				.param_width		(640),
				.param_height		(480),
				.param_awlen		(0), // (7),
				
				
				.monitor_addr		(),
				.monitor_stride		(),
				.monitor_width		(),
				.monitor_height		(),
				.monitor_awlen		(),
				
				.m_axi4_awid		(axi4_awid),
				.m_axi4_awaddr		(axi4_awaddr),
				.m_axi4_awburst		(axi4_awburst),
				.m_axi4_awcache		(axi4_awcache),
				.m_axi4_awlen		(axi4_awlen),
				.m_axi4_awlock		(axi4_awlock),
				.m_axi4_awprot		(axi4_awprot),
				.m_axi4_awqos		(axi4_awqos),
				.m_axi4_awregion	(axi4_awregion),
				.m_axi4_awsize		(axi4_awsize),
				.m_axi4_awvalid		(axi4_awvalid),
				.m_axi4_awready		(axi4_awready),
				.m_axi4_wstrb		(axi4_wstrb),
				.m_axi4_wdata		(axi4_wdata),
				.m_axi4_wlast		(axi4_wlast),
				.m_axi4_wvalid		(axi4_wvalid),
				.m_axi4_wready		(axi4_wready),
				.m_axi4_bid			(axi4_bid),
				.m_axi4_bresp		(axi4_bresp),
				.m_axi4_bvalid		(axi4_bvalid),
				.m_axi4_bready		(axi4_bready),
				
				.s_axi4s_tuser		(s_axi4s_tuser),
				.s_axi4s_tlast		(s_axi4s_tlast),
				.s_axi4s_tdata		(s_axi4s_tdata),
				.s_axi4s_tvalid		(s_axi4s_tvalid & ~s_axi4s_busy),
				.s_axi4s_tready		(s_axi4s_tready)
			);
	
	
	
	model_axi4_slave
			#(
				.AXI_ID_WIDTH		(AXI4_ID_WIDTH),
				.AXI_DATA_SIZE		(2),				// log2(n/8)  0:8bit, 1:16bit, 2:32bit, 3:64bit, ...
				.AXI_ADDR_WIDTH		(AXI4_ADDR_WIDTH),
				.AXI_QOS_WIDTH		(AXI4_QOS_WIDTH),
				.AXI_LEN_WIDTH		(AXI4_LEN_WIDTH),
				.MEM_SIZE			(4096)
			)
		i_model_axi4_slave
			(
				.aresetn			(~reset),
				.aclk				(clk),
				
				.s_axi4_awid		(axi4_awid),
				.s_axi4_awaddr		(axi4_awaddr),
				.s_axi4_awlen		(axi4_awlen),
				.s_axi4_awsize		(axi4_awsize),
				.s_axi4_awburst		(axi4_awburst),
				.s_axi4_awlock		(axi4_awlock),
				.s_axi4_awcache		(axi4_awcache),
				.s_axi4_awprot		(axi4_awprot),
				.s_axi4_awqos		(axi4_awqos),
				.s_axi4_awvalid		(axi4_awvalid),
				.s_axi4_awready		(axi4_awready),
				.s_axi4_wdata		(axi4_wdata),
				.s_axi4_wstrb		(axi4_wstrb),
				.s_axi4_wlast		(axi4_wlast),
				.s_axi4_wvalid		(axi4_wvalid),
				.s_axi4_wready		(axi4_wready),
				.s_axi4_bid			(axi4_bid),
				.s_axi4_bresp		(axi4_bresp),
				.s_axi4_bvalid		(axi4_bvalid),
				.s_axi4_bready		(axi4_bready),
				
				.s_axi4_arid		(axi4_arid),
				.s_axi4_araddr		(axi4_araddr),
				.s_axi4_arlen		(axi4_arlen),
				.s_axi4_arsize		(axi4_arsize),
				.s_axi4_arburst		(axi4_arburst),
				.s_axi4_arlock		(axi4_arlock),
				.s_axi4_arcache		(axi4_arcache),
				.s_axi4_arprot		(axi4_arprot),
				.s_axi4_arqos		(axi4_arqos),
				.s_axi4_arvalid		(axi4_arvalid),
				.s_axi4_arready		(axi4_arready),
				
				.s_axi4_rid			(axi4_rid),
				.s_axi4_rdata		(axi4_rdata),
				.s_axi4_rresp		(axi4_rresp),
				.s_axi4_rlast		(axi4_rlast),
				.s_axi4_rvalid		(axi4_rvalid),
				.s_axi4_rready		(axi4_rready)
			);

endmodule


`default_nettype wire


// end of file
